// ------------------------------------------------------
//-------------------- �������� ����� -------------------
// ------------------------------------------------------
parameter int BIT_RATE = 115200;    // �������� ������ � ���/�
parameter int BIT_PER_WORD = 8;     // ����� ��� � ����� ����� ������
parameter int PARITY_BIT = 1;       // ��� ���������: 0 - none, 1 - odd, 2 - even
parameter int STOP_BITS_NUM = 1;    // ����� ����-���: 1 ��� 2
