// ------------------------------------------------------
//-------------------- тестовый набор -------------------
// ------------------------------------------------------
parameter int BIT_RATE = 57600;     // скорость данных в бит/с
parameter int BIT_PER_WORD = 8;     // число бит в одном слове данных
parameter int PARITY_BIT = 0;       // бит четсности: 0 - none, 1 - odd, 2 - even
parameter int STOP_BITS_NUM = 1;    // число стоп-бит: 1 или 2
