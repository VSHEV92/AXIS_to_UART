// ------------------------------------------------------
//---------- ��������� ��������� ��������� --------------
// ------------------------------------------------------
parameter int CLK_FREQ = 100;              // �������� ������� � MHz  
parameter int RESET_DEASSERT_DELAY = 100;  // ����� ������ ������� ������ ns
parameter int DATA_WORDS_NUMB = 100;      // ����� ������������ ����
parameter int PARITY_ERR_PROB = 7;         // ������ � ������������ ����� � ���������

parameter int DATA_MIN_DELAY = 5*10e4;      // ������������ �������� ����� ��������� ������
parameter int DATA_MAX_DELAY = 10e5;      // ������������ �������� ����� ��������� ������
